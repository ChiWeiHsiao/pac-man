`timescale 1ns / 1ps
module pacman(
    input  clk,
    input  reset,//btn_s
	input  btn_n,
	input  btn_e,
	input  btn_w,
	input ROT_A,
	input ROT_B,
	input ROT_CENTER,
	input SW0,
	input SW1,
	input SW2,
	input SW3,
	output reg [7:0]led,
    // VGA specific I/O ports
    output HSYNC,
    output VSYNC,
    output VGA_RED,
    output VGA_GREEN,
    output VGA_BLUE
    );
wire rotary_event,rotary_right;

wire pixel_tick;    // when pixel tick is 1, we must update the RGB value
                    // based for the new coordinate (pixel_x, pixel_y)

wire [9:0] pixel_x; // x coordinate of the next pixel (between 0 ~ 639) 
wire [9:0] pixel_y; // y coordinate of the next pixel (between 0 ~ 479)

reg [2:0] rgb_reg;  // RGB value for the current pixel
reg [2:0] rgb_next; // RGB value for the next pixel

// Application-specific VGA signals
wire [2:0] current_rgb; // RGB values for the frame display application.
                        // In this demo, the value is generated by
                        // a video pattern generator:
                        //      video_pattern(id, x, y, current_rgb),
                        // where the input is the current scan coordinate (x, y),
                        // and the output is the RGB value of the video pattern
                        // 'id' at pixel (x, y).
// Declare system variables
wire [2:0]  btn_level, btn_pressed;
reg  [2:0]  prev_btn_level;

debounce btn_db0(
  .clk(clk),
  .btn_input(btn_n),
  .btn_output(btn_level[0])
  );

debounce btn_db1(
  .clk(clk),
  .btn_input(btn_e),
  .btn_output(btn_level[1])
  );
 
debounce btn_db2(
  .clk(clk),
  .btn_input(btn_w),
  .btn_output(btn_level[2])
  );
// instiantiate a VGA sync signal generator
vga_sync vs0(
  .clk(clk), .reset(reset), .oHS(HSYNC), .oVS(VSYNC),
  .visible(video_on), .p_tick(pixel_tick),
  .pixel_x(pixel_x), .pixel_y(pixel_y)
  );
  
Rotation_direction rotate(
    .CLK(clk),
    .ROT_A(ROT_A),
		.ROT_B(ROT_B),
		.rotary_event(rotary_event),
		.rotary_right(rotary_right)
    );

// Button click controller
always @(posedge clk) begin
  if (reset)
    prev_btn_level <= 3'b111;
  else
    prev_btn_level <= btn_level;
end

assign btn_pressed = (btn_level & ~prev_btn_level);

// VGA color pixel generator
assign {VGA_RED, VGA_GREEN, VGA_BLUE} = rgb_reg;

always @(posedge clk) begin
  if (pixel_tick)
    rgb_reg <= rgb_next;
  else
    rgb_reg <= rgb_reg;
end

always @(*) begin
  if (~video_on)
    rgb_next = 3'b000; // synchronization period, no need to set RGB values
  else
    rgb_next = current_rgb; // RGB value at (pixel_x, pixel_y)
end

//rotary
reg [9:0] rotary;
always@(posedge clk)begin
	if(reset) rotary<=0;
	else if(rotary_event && rotary_right && rotary < 60)//(640-16-32)/10
		rotary <= rotary+1;//讓count跑完一次週期中，亮的時間比例變長
	else if(rotary_event && !rotary_right && rotary>0)
		rotary <= rotary-1;
	else rotary <= rotary;
end
//----------------------------------------------------------------------------------------------------------------------
//控制11個tp下落的時間
reg [20:0] tp_time;
reg [20:0]tp_cnt;//除頻
reg tp_start_to_fall;
always@(posedge clk)begin
	if(reset) tp_start_to_fall<=0;
	else if(ROT_CENTER)tp_start_to_fall<=1;
end
always@(posedge clk)begin
	if(reset)begin
		tp_cnt<=0;
		tp_time<=0; end
	else if(tp_start_to_fall) begin
		if(SW3) begin tp_cnt <= tp_cnt; tp_time <= tp_time; end// pause
		else if(tp_cnt == 500000)begin//設成500000->0.01sec
			tp_cnt<=0;
			tp_time <= tp_time+1;end
		else 
			tp_cnt <= tp_cnt + 1;
	end
end
// 畫gp 嘴巴會動的小精靈
wire gp_pattern[0:31][0:31];
`include "gp_pattern.dat"
wire gp_pattern2[0:31][0:31];
`include "gp_pattern2.dat"
wire gp_on;
reg [9:0]gp_x, gp_y;//gp左上的參考點
reg mouth;
reg [30:0]mouth_cnt;
always@(posedge clk) begin
	if(reset)begin mouth<=0; mouth_cnt<=0;end
	else 
		if(mouth_cnt == 5000000)begin//除頻 5000000->0.1sec
			mouth_cnt<=0;
			mouth<=!mouth;end
		else mouth_cnt <= mouth_cnt + 1;
end

assign gp_on = mouth ?
				((pixel_x>=gp_x && pixel_x<=gp_x+32) && (pixel_y>=gp_y && pixel_y<=gp_y+32) && gp_pattern[pixel_x-gp_x][pixel_y-gp_y]) : 
				((pixel_x>=gp_x && pixel_x<=gp_x+32) && (pixel_y>=gp_y && pixel_y<=gp_y+32) && gp_pattern2[pixel_x-gp_x][pixel_y-gp_y]);


always@(posedge clk) begin
	gp_x<=0 + (rotary*10); //*10 改改改 <<3
	gp_y<=480-32;
end
//畫circle
wire circle_pattern[0:19][0:19];
`include "circle_pattern.dat"
//畫triangle
wire triangle_pattern[0:19][0:19];
`include "triangle_pattern.dat"
//畫square
wire square_pattern[0:19][0:19];
`include "square_pattern.dat"

//reg [9:0]bullet_x, bullet_y;
reg [9:0] get_x;
reg [9:0] cnt_x;//random position of TP (0~640-20)
always@(posedge clk)begin
	if(reset)begin
		cnt_x<=0;
		get_x<=0; end
	else begin
		if(ROT_CENTER) get_x <= cnt_x;
	
		if(cnt_x == 640-20) cnt_x <= 0;
		else cnt_x <= cnt_x+1;
	end
end

//tp t0~10
`include "c0.dat"//1 
`include "t1.dat"//100
`include "c2.dat"//130
`include "s3.dat"//200
`include "t4.dat"//t4 280 
`include "t5.dat"//t5 355 
`include "s6.dat"//s6 490
`include "c7.dat"//c7 570 
`include "s8.dat"//s8 650
`include "s9.dat"//s9 830
`include "t10.dat"//t10 900 

//畫status board 剩下幾個tp要掉落
`include "zero.dat"
`include "one.dat"
`include "two.dat"
`include "three.dat"
`include "four.dat"
`include "five.dat"
`include "six.dat"
`include "seven.dat"
`include "eight.dat"
`include "nine.dat"
`include "ten.dat"
`include "eleven.dat"
reg [4:0]remain_tp;
assign zero_on=(remain_tp==0 && (pixel_x>=550 && pixel_x<590) && (pixel_y>=50 && pixel_y<90) && zero[pixel_x-550][pixel_y-50]);
assign one_on=(remain_tp==1 && (pixel_x>=550 && pixel_x<590) && (pixel_y>=50 && pixel_y<90) && one[pixel_x-550][pixel_y-50]);
assign two_on=(remain_tp==2 && (pixel_x>=550 && pixel_x<590) && (pixel_y>=50 && pixel_y<90) && two[pixel_x-550][pixel_y-50]);
assign three_on=(remain_tp==3 && (pixel_x>=550 && pixel_x<590) && (pixel_y>=50 && pixel_y<90) && three[pixel_x-550][pixel_y-50]);
assign four_on=(remain_tp==4 && (pixel_x>=550 && pixel_x<590) && (pixel_y>=50 && pixel_y<90) && four[pixel_x-550][pixel_y-50]);
assign five_on=(remain_tp==5 && (pixel_x>=550 && pixel_x<590) && (pixel_y>=50 && pixel_y<90) && five[pixel_x-550][pixel_y-50]);
assign six_on=(remain_tp==6 && (pixel_x>=550 && pixel_x<590) && (pixel_y>=50 && pixel_y<90) && six[pixel_x-550][pixel_y-50]);
assign seven_on=(remain_tp==7 && (pixel_x>=550 && pixel_x<590) && (pixel_y>=50 && pixel_y<90) && seven[pixel_x-550][pixel_y-50]);
assign eight_on=(remain_tp==8 && (pixel_x>=550 && pixel_x<590) && (pixel_y>=50 && pixel_y<90) && eight[pixel_x-550][pixel_y-50]);
assign nine_on=(remain_tp==9 && (pixel_x>=550 && pixel_x<590) && (pixel_y>=50 && pixel_y<90) && nine[pixel_x-550][pixel_y-50]);
assign ten_on=(remain_tp==10 && (pixel_x>=550 && pixel_x<590) && (pixel_y>=50 && pixel_y<90) && ten[pixel_x-550][pixel_y-50]);
assign eleven_on=(remain_tp==11 && (pixel_x>=550 && pixel_x<590) && (pixel_y>=50 && pixel_y<90) && eleven[pixel_x-550][pixel_y-50]);

wire status_on;//40*40
assign status_on = ((pixel_x>=550 && pixel_x<=590) && (pixel_y>=50 && pixel_y<=90))?1:0;
always@(posedge clk) begin //算剩下的數量
	if(reset)begin remain_tp<=11;end
	else begin
		if(tp_time==1||tp_time==200||tp_time==250||tp_time==350||tp_time==400||tp_time==550||tp_time==600||tp_time==750||tp_time==870||tp_time==950||tp_time==1100)
			remain_tp <= remain_tp-1;
	end
end
//判斷gp是否有吃到tp
reg [4:0] total_got;
reg [4:0] circle_got;
reg [4:0] square_got;
reg [4:0] triangle_got;
always@(posedge clk)begin
	if(reset) begin
		total_got<=0; circle_got<=0; square_got<=0; triangle_got<=0; end
	else begin
		if((c0_x>=gp_x-20 && c0_x<=gp_x+32) && gp_y==c0_y)begin circle_got<= circle_got+1; total_got <= total_got+1;end
		if((t1_x>=gp_x-20 && t1_x<=gp_x+32) && gp_y==t1_y)begin triangle_got<= triangle_got+1; total_got<= total_got+1;end
		if((c2_x>=gp_x-20 && c2_x<=gp_x+32) && gp_y==c2_y)begin circle_got<= circle_got+1; total_got<= total_got+1;end
		if((s3_x>=gp_x-20 && s3_x<=gp_x+32) && gp_y==s3_y)begin square_got<= square_got+1; total_got<= total_got+1;end
		if((t4_x>=gp_x-20 && t4_x<=gp_x+32) && gp_y==t4_y)begin triangle_got<= triangle_got+1; total_got<= total_got+1;end
		if((t5_x>=gp_x-20 && t5_x<=gp_x+32) && gp_y==t5_y)begin triangle_got<= triangle_got+1; total_got<= total_got+1;end
		if((s6_x>=gp_x-20 && s6_x<=gp_x+32) && gp_y==s6_y)begin square_got<= square_got+1; total_got<= total_got+1;end
		if((c7_x>=gp_x-20 && c7_x<=gp_x+32) && gp_y==c7_y)begin circle_got<= circle_got+1; total_got<= total_got+1;end
		if((s8_x>=gp_x-20 && s8_x<=gp_x+32) && gp_y==s8_y)begin square_got<= square_got+1; total_got<= total_got+1;end
		if((s9_x>=gp_x-20 && s9_x<=gp_x+32) && gp_y==s9_y)begin square_got<= square_got+1; total_got<= total_got+1;end
		if((t10_x>=gp_x-20 && t10_x<=gp_x+32) && gp_y==t10_y)begin triangle_got<= triangle_got+1; total_got<= total_got+1;end
	end
end

//Final score board 分別顯示有幾個有幾個三角形圓形正方形 改改改
wire final_on;//40*40
assign final_on = (tp_time>=1100+480 && (pixel_x>=100 && pixel_x<=400) && (pixel_y>=150 && pixel_y<=400) && !circle_pattern[pixel_x-150][pixel_y-200] && !triangle_pattern[pixel_x-150][pixel_y-260] && !square_pattern[pixel_x-150][pixel_y-310]);
wire score_c_on;//40*40 (200,180)
assign score_c_on = (tp_time>=1100+480 && circle_got==0)? (pixel_x>=200 && pixel_x<=240 && pixel_y>=180 && pixel_y<=220 && zero[pixel_x-200][pixel_y-180]):
					(tp_time>=1100+480 && circle_got==1)? (pixel_x>=200 && pixel_x<=240 && pixel_y>=180 && pixel_y<=220 && one[pixel_x-200][pixel_y-180]):
					(tp_time>=1100+480 && circle_got==2)? (pixel_x>=200 && pixel_x<=240 && pixel_y>=180 && pixel_y<=220 && two[pixel_x-200][pixel_y-180]):
					(tp_time>=1100+480 && circle_got==3)? (pixel_x>=200 && pixel_x<=240 && pixel_y>=180 && pixel_y<=220 && three[pixel_x-200][pixel_y-180]):
					(tp_time>=1100+480 && circle_got==4)? (pixel_x>=200 && pixel_x<=240 && pixel_y>=180 && pixel_y<=220 && four[pixel_x-200][pixel_y-180]):
					0;

wire score_t_on;//40*40 (200,240)
assign score_t_on = (tp_time>=1100+480 && triangle_got==0)? (pixel_x>=200 && pixel_x<=240 && pixel_y>=240 && pixel_y<=280 && zero[pixel_x-200][pixel_y-240]):
					(tp_time>=1100+480 && triangle_got==1)? (pixel_x>=200 && pixel_x<=240 && pixel_y>=240 && pixel_y<=280 && one[pixel_x-200][pixel_y-240]):
					(tp_time>=1100+480 && triangle_got==2)? (pixel_x>=200 && pixel_x<=240 && pixel_y>=240 && pixel_y<=280 && two[pixel_x-200][pixel_y-240]):
					(tp_time>=1100+480 && triangle_got==3)? (pixel_x>=200 && pixel_x<=240 && pixel_y>=240 && pixel_y<=280 && three[pixel_x-200][pixel_y-240]):
					(tp_time>=1100+480 && triangle_got==4)? (pixel_x>=200 && pixel_x<=240 && pixel_y>=240 && pixel_y<=280 && four[pixel_x-200][pixel_y-240]):
					0;
					
wire score_s_on;//40*40 (200,300)
assign score_s_on = (tp_time>=1100+480 && square_got==0)? (pixel_x>=200 && pixel_x<=240 && pixel_y>=300 && pixel_y<=340 && zero[pixel_x-200][pixel_y-300]):
					(tp_time>=1100+480 && square_got==1)? (pixel_x>=200 && pixel_x<=240 && pixel_y>=300 && pixel_y<=340 && one[pixel_x-200][pixel_y-300]):
					(tp_time>=1100+480 && square_got==2)? (pixel_x>=200 && pixel_x<=240 && pixel_y>=300 && pixel_y<=340 && two[pixel_x-200][pixel_y-300]):
					(tp_time>=1100+480 && square_got==3)? (pixel_x>=200 && pixel_x<=240 && pixel_y>=300 && pixel_y<=340 && three[pixel_x-200][pixel_y-300]):
					(tp_time>=1100+480 && square_got==4)? (pixel_x>=200 && pixel_x<=240 && pixel_y>=300 && pixel_y<=340 && four[pixel_x-200][pixel_y-300]):
					0;
//switch change gp color
//0=red; 1=green; 2=blue; 0+1=plain blue; 0+2=pink; 1+2=yello; all=white;
reg r_on, g_on, b_on;//color
always@(posedge clk)begin
	if(SW2)begin//gp 0+1+2
		r_on <= score_t_on || score_s_on || score_c_on || gp_on || c2_on || s3_on || t5_on || s9_on || t4_on || c7_on || s8_on || bullet_on;
		g_on <= final_on||gp_on || c0_on || t10_on || s3_on || t4_on || c7_on || zero_on || one_on || two_on || three_on || three_on || four_on || five_on || six_on || seven_on || eight_on || nine_on || ten_on || eleven_on;
		b_on <= gp_on || status_on || t1_on || s6_on || t5_on || s9_on || t4_on || c7_on ;end
	else if(SW1)begin//gp 0+2
		r_on <= score_t_on || score_s_on || score_c_on || gp_on || c2_on || s3_on || t5_on || s9_on || t4_on || c7_on || s8_on || bullet_on;
		g_on <= final_on||c0_on || t10_on || s3_on || t4_on || c7_on || zero_on ||  one_on || two_on || three_on || three_on || four_on || five_on || six_on || seven_on || eight_on || nine_on || ten_on || eleven_on;
		b_on <= gp_on || status_on || t1_on || s6_on || t5_on || s9_on || t4_on || c7_on ;end
	else if(SW0)begin//gp 0+1
		r_on <= score_t_on || score_s_on || score_c_on || gp_on || c2_on || s3_on || t5_on || s9_on || t4_on || c7_on || s8_on || bullet_on;
		g_on <= final_on||gp_on || c0_on || t10_on || s3_on || t4_on || c7_on || zero_on ||  one_on || two_on || three_on || three_on || four_on || five_on || six_on || seven_on || eight_on || nine_on || ten_on || eleven_on;
		b_on <= t1_on || status_on || s6_on || t5_on || s9_on || t4_on || c7_on ;end
	else begin//yellow 1+2
		r_on <= score_t_on || score_s_on || score_c_on || c2_on || s3_on || t5_on || s9_on || t4_on || c7_on || s8_on || bullet_on;
		g_on <= final_on||gp_on || c0_on || t10_on || s3_on || t4_on || c7_on || zero_on ||  one_on || two_on || three_on || three_on || four_on || five_on || six_on || seven_on || eight_on || nine_on || ten_on || eleven_on;
		b_on <= gp_on || status_on || t1_on || s6_on || t5_on || s9_on || t4_on || c7_on ;end
end
//score_t_on || score_s_on || score_c_on || 
//current_rgb 顯示 xx_on 
assign current_rgb[0] = r_on;
assign current_rgb[1] = g_on;
assign current_rgb[2] = b_on;

//led顯示得分
always@(posedge clk)begin
	if(reset) led <= 8'd0;
	else led <= total_got;//total_got
end

endmodule
