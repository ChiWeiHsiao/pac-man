`timescale 1ns / 1ps
module final(
    input  clk,
    input  reset,//btn_s
	 input  btn_n,
	 input  btn_e,
	 input  btn_w,

    // VGA specific I/O ports
    output HSYNC,
    output VSYNC,
    output VGA_RED,
    output VGA_GREEN,
    output VGA_BLUE
    );

// general VGA control signals
//wire video_on;      // when video_on is 0, the VGA controller is sending
                    // synchronization signals to the display device.

wire pixel_tick;    // when pixel tick is 1, we must update the RGB value
                    // based for the new coordinate (pixel_x, pixel_y)

wire [9:0] pixel_x; // x coordinate of the next pixel (between 0 ~ 639) 
wire [9:0] pixel_y; // y coordinate of the next pixel (between 0 ~ 479)

/* �e�� x^2+y^<r^
reg [9:0] centerx;//��ߪ�x�y��
reg [9:0] centery;//��ߪ�y�y��
wire [19:0] xsq;
wire [19:0] ysq;
assign xsq = (pixel_x-centerx)*(pixel_x-centerx);
assign ysq = (pixel_y-centery)*(pixel_y-centery);*/

reg [2:0] rgb_reg;  // RGB value for the current pixel
reg [2:0] rgb_next; // RGB value for the next pixel

// Application-specific VGA signals
reg [2:0] current_rgb; // RGB values for the frame display application.
                        // In this demo, the value is generated by
                        // a video pattern generator:
                        //      video_pattern(id, x, y, current_rgb),
                        // where the input is the current scan coordinate (x, y),
                        // and the output is the RGB value of the video pattern
                        // 'id' at pixel (x, y).
								
reg  [2:0] pattern_id;// circle, triangle, square

// Declare system variables
wire [2:0]  btn_level, btn_pressed;
reg  [2:0]  prev_btn_level;
reg  [8:0] sd_counter;

debounce btn_db0(
  .clk(clk),
  .btn_input(btn_n),
  .btn_output(btn_level[0])
  );

debounce btn_db1(
  .clk(clk),
  .btn_input(btn_e),
  .btn_output(btn_level[1])
  );
 
debounce btn_db2(
  .clk(clk),
  .btn_input(btn_w),
  .btn_output(btn_level[2])
  );
// instiantiate a VGA sync signal generator
vga_sync vs0(
  .clk(clk), .reset(reset), .oHS(HSYNC), .oVS(VSYNC),
  .visible(video_on), .p_tick(pixel_tick),
  .pixel_x(pixel_x), .pixel_y(pixel_y)
  );
clk_divider#(100) clk_divider0(
    .clk(clk),
    .reset(reset),
    .clk_out(clk_500k)
  );

// Button click controller
always @(posedge clk) begin
  if (reset)
    prev_btn_level <= 3'b111;
  else
    prev_btn_level <= btn_level;
end

assign btn_pressed = (btn_level & ~prev_btn_level);

// VGA color pixel generator
assign {VGA_RED, VGA_GREEN, VGA_BLUE} = rgb_reg;

always @(posedge clk) begin
  if (pixel_tick)
    rgb_reg <= rgb_next;
  else
    rgb_reg <= rgb_reg;
end

always @(*) begin
  if (~video_on)
    rgb_next = 3'b000; // synchronization period, no need to set RGB values
  else
    rgb_next = current_rgb; // RGB value at (pixel_x, pixel_y)
end
//----------------------------------------------------------------------------------------------------------------------
// �egp array
wire gp_pattern[0:31][0:31];
`include "gp_pattern.dat"
wire gp_on;
reg [9:0]gp_x, gp_y;
assign gp_on = ((pixel_x>=gp_x && pixel_x<=gp_x+32) && (pixel_y>=gp_y && pixel_y<=gp_y+32) && gp_pattern[pixel_x-gp_x][pixel_y-gp_y])?1:0;
always@(posedge clk) begin
  gp_x<=100; gp_y<=100;//gp���W���Ѧ��I
end
//�ecircle
wire circle_pattern[0:19][0:19];
`include "circle_pattern.dat"
wire circle_on;
reg [9:0]circle_x, circle_y;
assign circle_on = ((pixel_x>=circle_x && pixel_x<=circle_x+20) && (pixel_y>=circle_y && pixel_y<=circle_y+20) && circle_pattern[pixel_x-circle_x][pixel_y-circle_y])?1:0;
always@(posedge clk) begin
  circle_x<=150; circle_y<=150;//circle���W���Ѧ��I
end
//�etriangle
wire triangle_pattern[0:19][0:19];
`include "triangle_pattern.dat"
wire triangle_on;
reg [9:0]triangle_x, triangle_y;
assign triangle_on = ((pixel_x>=triangle_x && pixel_x<=triangle_x+20) && (pixel_y>=triangle_y && pixel_y<=triangle_y+20) && triangle_pattern[pixel_x-triangle_x][pixel_y-triangle_y])?1:0;
always@(posedge clk) begin
  triangle_x<=150; triangle_y<=100;//circle���W���Ѧ��I
end
//�esquare
wire square_pattern[0:19][0:19];
`include "square_pattern.dat"
wire square_on;
reg [9:0]square_x, square_y;
assign square_on = ((pixel_x>=square_x && pixel_x<=square_x+20) && (pixel_y>=square_y && pixel_y<=square_y+20) && square_pattern[pixel_x-square_x][pixel_y-square_y])?1:0;
always@(posedge clk) begin
  square_x<=60; square_y<=200;//circle���W���Ѧ��I
end

//pixel_x,y  try
always @(posedge clk) begin
	current_rgb[0] <=gp_on || circle_on || triangle_on || square_on;
	current_rgb[2] <=gp_on || circle_on || triangle_on || square_on;
	/*
	if ( (pixel_x>=400 && pixel_x<=405) && (pixel_y>=100 && pixel_y<=150)) current_rgb <= 3'b010;//line
	else if() current_rgb <= 3'b111;//gp
	else if( (xsq+ysq)<1024) current_rgb <= 3'b111;//circle
	else current_rgb <= 3'b000;//background
	*/
end

endmodule
